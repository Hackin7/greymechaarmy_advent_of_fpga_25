module coprocessor(
    input clk, 
    input rst, 
    input data_valid
);
endmodule